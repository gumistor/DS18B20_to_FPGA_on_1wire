`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Asynchronous driver
//////////////////////////////////////////////////////////////////////////////////
module ram (reset, din, write_en, waddr, wclk, raddr, rclk, dout);//512x8
 parameter addr_width = 9;
 parameter data_width = 8;
 input [addr_width-1:0] waddr, raddr;
 input [data_width-1:0] din;
 input reset;
 input write_en, wclk, rclk;
 output reg [data_width-1:0] dout;
 reg [data_width-1:0] mem [(1<<addr_width)-1:0];
 
 initial $readmemh("C:\\Users\\Krzysztof\\Documents\\fpga_temperature_sensor\\memory.dat", mem);
 
 always @(posedge wclk) // Write memory.
 begin
	if (write_en)
		mem[waddr] <= din; // Using write address bus.
end

always @(posedge rclk) // Read memory.
if(reset) dout <= 8'h0;
else
	begin
		dout <= mem[raddr]; // Using read address bus.
	end
 /*
parameter INIT_0 = 
256'h54797369613a2a2030303A30303A30302B3030302C30303030DF432020202020;
parameter INIT_1 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_2 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_3 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_4 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_5 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_6 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_7 = 
256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_9 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_A = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_B = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_C = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_D = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_E = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
parameter INIT_F = 
256'h0000000000000000000000000000000000000000000000000000000000000000;
 */
endmodule
/*
defparam ram512x8_inst.INIT_0 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_1 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_2 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_3 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_4 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_5 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_6 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_7 = 
256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram512x8_inst.INIT_8 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_9 = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_A = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_B = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_C = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_D = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_E = 
256'h0000000000000000000000000000000000000000000000000000000000000000; 
defparam ram512x8_inst.INIT_F = 
256'h0000000000000000000000000000000000000000000000000000000000000000;
*/